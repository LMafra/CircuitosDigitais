library verilog;
use verilog.vl_types.all;
entity coder_vlg_sample_tst is
    port(
        S1              : in     vl_logic;
        S2              : in     vl_logic;
        S3              : in     vl_logic;
        S4              : in     vl_logic;
        S5              : in     vl_logic;
        S6              : in     vl_logic;
        S7              : in     vl_logic;
        S8              : in     vl_logic;
        S9              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end coder_vlg_sample_tst;
