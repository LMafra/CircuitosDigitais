library verilog;
use verilog.vl_types.all;
entity coder_vlg_vec_tst is
end coder_vlg_vec_tst;
